LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY bcd_7segment IS
	PORT (
		bcd_in : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		seven_segment_out : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		seven_segment_out1 : OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
	);
END bcd_7segment;

ARCHITECTURE Behavioral OF bcd_7segment IS
BEGIN
	PROCESS (bcd_in)
	BEGIN
		CASE bcd_in IS
			WHEN "00000000" => -- x0
				seven_segment_out <= NOT "0111111";
				seven_segment_out1 <= NOT "0000000";
			WHEN "00000001" => --x1
				seven_segment_out <= NOT "0000110";
				seven_segment_out1 <= NOT "0000000";
			WHEN "00000010" => --x2
				seven_segment_out <= NOT "1011011";
				seven_segment_out1 <= NOT "0000000";
			WHEN "00000011" => --x3
				seven_segment_out <= NOT "1001111";
				seven_segment_out1 <= NOT "0000000";
			WHEN "00000100" => --x4
				seven_segment_out <= NOT "1100110";
				seven_segment_out1 <= NOT "0000000";
			WHEN "00000101" => --x5
				seven_segment_out <= NOT "1101101";
				seven_segment_out1 <= NOT "0000000";
			WHEN "00000110" => --x6
				seven_segment_out <= NOT "1111101";
				seven_segment_out1 <= NOT "0000000";
			WHEN "00000111" => --x7
				seven_segment_out <= NOT "0000111";
				seven_segment_out1 <= NOT "0000000";
			WHEN "00001000" => --x8
				seven_segment_out <= NOT "1111111";
				seven_segment_out1 <= NOT "0000000";
			WHEN "00001001" => --x9
				seven_segment_out <= NOT "1100111";
				seven_segment_out1 <= NOT "0000000";
			WHEN "00001010" => -- 10
				seven_segment_out <= NOT "0111111";
				seven_segment_out1 <= NOT "0000110";
			WHEN "00001011" => --11
				seven_segment_out <= NOT "0000110";
				seven_segment_out1 <= NOT "0000110";
			WHEN "00001100" => --12
				seven_segment_out <= NOT "1011011";
				seven_segment_out1 <= NOT "0000110";
			WHEN "00001101" => --13
				seven_segment_out <= NOT "1001111";
				seven_segment_out1 <= NOT "0000110";
			WHEN "00001110" => --14
				seven_segment_out <= NOT "1100110";
				seven_segment_out1 <= NOT "0000110";
			WHEN "00001111" => --15
				seven_segment_out <= NOT "1101101";
				seven_segment_out1 <= NOT "0000110";
			WHEN "00010000" => -- 16
				seven_segment_out <= NOT "1111101";
				seven_segment_out1 <= NOT "0000110";
			WHEN "00010001" => -- 17
				seven_segment_out <= NOT "0000111";
				seven_segment_out1 <= NOT "0000110";
			WHEN "00010010" => -- 18
				seven_segment_out <= NOT "1111111";
				seven_segment_out1 <= NOT "0000110";
			WHEN "00010011" => -- 19
				seven_segment_out <= NOT "1100111";
				seven_segment_out1 <= NOT "0000110";
			WHEN "00010100" => -- 20
				seven_segment_out <= NOT "0111111";
				seven_segment_out1 <= NOT "1011011";
			WHEN "00010101" => -- 21
				seven_segment_out <= NOT "0000110";
				seven_segment_out1 <= NOT "1011011";
			WHEN "00010110" => -- 22
				seven_segment_out <= NOT "1011011";
				seven_segment_out1 <= NOT "1011011";
			WHEN "00010111" => -- 23
				seven_segment_out <= NOT "1001111";
				seven_segment_out1 <= NOT "1011011";
			WHEN "00011000" => -- 24
				seven_segment_out <= NOT "1100110";
				seven_segment_out1 <= NOT "1011011";
			WHEN "00011001" => -- 25
				seven_segment_out <= NOT "1101101";
				seven_segment_out1 <= NOT "1011011";
			WHEN "00011010" => -- 26
				seven_segment_out <= NOT "1111101";
				seven_segment_out1 <= NOT "1011011";
			WHEN "00011011" => -- 27
				seven_segment_out <= NOT "0000111";
				seven_segment_out1 <= NOT "1011011";
			WHEN "00011100" => -- 28
				seven_segment_out <= NOT "1111111";
				seven_segment_out1 <= NOT "1011011";
			WHEN "00011101" => -- 29
				seven_segment_out <= NOT "1100111";
				seven_segment_out1 <= NOT "1011011";
			WHEN "00011110" => -- 30
				seven_segment_out <= NOT "0111111";
				seven_segment_out1 <= NOT "1001111";
			WHEN "00011111" => -- 31
				seven_segment_out <= NOT "0000110";
				seven_segment_out1 <= NOT "1001111";
			WHEN "00100000" => -- 32
				seven_segment_out <= NOT "1011011";
				seven_segment_out1 <= NOT "1001111";
			WHEN "00100001" => -- 33
				seven_segment_out <= NOT "1001111";
				seven_segment_out1 <= NOT "1001111";
			WHEN "00100010" => -- 34
				seven_segment_out <= NOT "1100110";
				seven_segment_out1 <= NOT "1001111";
			WHEN "00100011" => -- 35
				seven_segment_out <= NOT "1101101";
				seven_segment_out1 <= NOT "1001111";
			WHEN "00100100" => -- 36
				seven_segment_out <= NOT "1111101";
				seven_segment_out1 <= NOT "1001111";
			WHEN "00100101" => -- 37
				seven_segment_out <= NOT "0000111";
				seven_segment_out1 <= NOT "1001111";
			WHEN "00100110" => -- 38
				seven_segment_out <= NOT "1111111";
				seven_segment_out1 <= NOT "1001111";
			WHEN "00100111" => -- 39
				seven_segment_out <= NOT "1100111";
				seven_segment_out1 <= NOT "1001111";
			WHEN "00101000" => -- 40
				seven_segment_out <= NOT "0111111";
				seven_segment_out1 <= NOT "1100110";
			WHEN "00101001" => -- 41
				seven_segment_out <= NOT "0000110";
				seven_segment_out1 <= NOT "1100110";
			WHEN "00101010" => -- 42
				seven_segment_out <= NOT "1011011";
				seven_segment_out1 <= NOT "1100110";
			WHEN "00101011" => -- 43
				seven_segment_out <= NOT "1001111";
				seven_segment_out1 <= NOT "1100110";
			WHEN "00101100" => -- 44
				seven_segment_out <= NOT "1100110";
				seven_segment_out1 <= NOT "1100110";
			WHEN "00101101" => -- 45
				seven_segment_out <= NOT "1101101";
				seven_segment_out1 <= NOT "1100110";
			WHEN "00101110" => -- 46
				seven_segment_out <= NOT "1111101";
				seven_segment_out1 <= NOT "1100110";
			WHEN "00101111" => -- 47
				seven_segment_out <= NOT "0000111";
				seven_segment_out1 <= NOT "1100110";
			WHEN "00110000" => -- 48
				seven_segment_out <= NOT "1111111";
				seven_segment_out1 <= NOT "1100110";
			WHEN "00110001" => -- 49
				seven_segment_out <= NOT "1100111";
				seven_segment_out1 <= NOT "1100110";
			WHEN "00110010" => -- 50
				seven_segment_out <= NOT "0111111";
				seven_segment_out1 <= NOT "1101101";
			WHEN "00110011" => -- 51
				seven_segment_out <= NOT "0000110";
				seven_segment_out1 <= NOT "1101101";
			WHEN "00110100" => -- 52
				seven_segment_out <= NOT "1011011";
				seven_segment_out1 <= NOT "1101101";
			WHEN "00110101" => -- 53
				seven_segment_out <= NOT "1001111";
				seven_segment_out1 <= NOT "1101101";
			WHEN "00110110" => -- 54
				seven_segment_out <= NOT "1100110";
				seven_segment_out1 <= NOT "1101101";
			WHEN "00110111" => -- 55
				seven_segment_out <= NOT "1101101";
				seven_segment_out1 <= NOT "1101101";
			WHEN "00111000" => -- 56
				seven_segment_out <= NOT "1111101";
				seven_segment_out1 <= NOT "1101101";
			WHEN "00111001" => -- 57
				seven_segment_out <= NOT "0000111";
				seven_segment_out1 <= NOT "1101101";
			WHEN "0111010" => -- 58
				seven_segment_out <= NOT "1111111";
				seven_segment_out1 <= NOT "1101101";
			WHEN "00111011" => -- 59
				seven_segment_out <= NOT "1100111";
				seven_segment_out1 <= NOT "1101101";
			WHEN "00111100" => -- 60
				seven_segment_out <= NOT "0111111";
				seven_segment_out1 <= NOT "1111101";
			WHEN "00111101" => -- 61
				seven_segment_out <= NOT "0000110";
				seven_segment_out1 <= NOT "1111101";
			WHEN "00111110" => -- 62
				seven_segment_out <= NOT "1011011";
				seven_segment_out1 <= NOT "1111101";
			WHEN "00111111" => -- 63
				seven_segment_out <= NOT "1001111";
				seven_segment_out1 <= NOT "1111101";
 
			WHEN "01000000" => -- 64
				seven_segment_out <= NOT "1111110";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01000001" => -- 65
				seven_segment_out <= NOT "0110000";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01000010" => -- 66
				seven_segment_out <= NOT "1101101";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01000011" => -- 67
				seven_segment_out <= NOT "1111001";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01000100" => -- 68
				seven_segment_out <= NOT "1111111";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01000101" => -- 69
				seven_segment_out <= NOT "1110111";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01000110" => -- 70
				seven_segment_out <= NOT "1111011";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01000111" => -- 71
				seven_segment_out <= NOT "1111110";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01001000" => -- 72
				seven_segment_out <= NOT "0111001";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01001001" => -- 73
				seven_segment_out <= NOT "1011110";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01001010" => -- 74
				seven_segment_out <= NOT "1111100";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01001011" => -- 75
				seven_segment_out <= NOT "1111100";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01001100" => -- 76
				seven_segment_out <= NOT "0111000";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01001101" => -- 77
				seven_segment_out <= NOT "1111111";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01001110" => -- 78
				seven_segment_out <= NOT "1111000";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01001111" => -- 79
				seven_segment_out <= NOT "0111111";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01010000" => -- 80
				seven_segment_out <= NOT "1111111";
				seven_segment_out1 <= NOT "1111110"; 
			WHEN "01010001" => -- 81
				seven_segment_out <= NOT "1111001";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01010010" => -- 82
				seven_segment_out <= NOT "1110010";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01010011" => -- 83
				seven_segment_out <= NOT "1110110";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01010100" => -- 84
				seven_segment_out <= NOT "1111101";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01010101" => -- 85
				seven_segment_out <= NOT "1110111";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01010110" => -- 86
				seven_segment_out <= NOT "1111111";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01010111" => -- 87
				seven_segment_out <= NOT "1111001";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01011000" => -- 88
				seven_segment_out <= NOT "0111111";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01011001" => -- 89
				seven_segment_out <= NOT "1011111";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01011010" => -- 90
				seven_segment_out <= NOT "1111100";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01011011" => -- 91
				seven_segment_out <= NOT "1111110";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01011100" => -- 92
				seven_segment_out <= NOT "1111011";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01011101" => -- 93
				seven_segment_out <= NOT "0111001";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01011110" => -- 94
				seven_segment_out <= NOT "1101001";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01011111" => -- 95
				seven_segment_out <= NOT "1001111";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01100000" => -- 96
				seven_segment_out <= NOT "1111010";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01100001" => -- 97
				seven_segment_out <= NOT "1110000";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01100010" => -- 98
				seven_segment_out <= NOT "1001110";
				seven_segment_out1 <= NOT "1111110";
			WHEN "01100011" => -- 99
				seven_segment_out <= NOT "0001111";
				seven_segment_out1 <= NOT "1111110";
 
 
			WHEN OTHERS => 
				seven_segment_out <= NOT "1000000";
				seven_segment_out1 <= NOT "1000000";
		END CASE;
	END PROCESS;
END Behavioral;